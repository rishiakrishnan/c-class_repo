
/*
See LICENSE for details
This file has been generated by CSR-BOX - 1.7.0
Time of Generation: 2025-04-11 18:28:29.634185
*/

package csr_types ;
    `include "csrbox.defines"
    `include "Logger.bsv"


    typedef struct {
        Bit#(12) csr_address;
        Bit#(64) writedata;
        Bit#(2) funct3;
        Bit#(1) pc_1;
    } CSRReq deriving(Bits, FShow, Eq);

    typedef struct{
        Bool hit;
        Bit#(64)  data;
    `ifdef rtldump
        Bool csr_updated;
    `endif
    } CSRResponse deriving(Bits, Eq, FShow);

    typedef enum {Machine = 3, Hypervisor=2, Supervisor = 1, User = 0} Privilege_mode deriving(Bits, Eq, FShow);


    function Bit#(64) fn_csr_op (Bit#(64) writedata, Bit#(64) readdata, Bit#(2) op);
        if(op == 'd1)
    	    return writedata;
        else if(op == 'd2)
            return (writedata|readdata);
        else
            return (~writedata & readdata);
    endfunction
  
  function Reg#(Bit#(1)) extInterruptReg(Reg#(Bit#(1)) r1, Reg#(Bit#(1)) r2);
    return (interface Reg;
      method Bit#(1) _read = r1 | r2;
      method Action _write(Bit#(1) x);
        r1._write(x);
			endmethod
    endinterface);
  endfunction
  
endpackage 
