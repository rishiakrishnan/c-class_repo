
/*
See LICENSE for details
This file has been generated by CSR-BOX - 1.7.0
Time of Generation: 2025-04-11 18:28:29.636361
*/

package csrbox_grp1;
   
import Vector           :: *;
import FIFOF            :: * ;
import DReg             :: * ;
import UniqueWrappers   :: * ;
import ConcatReg        :: * ;
import GetPut           :: * ;
import Connectable      :: * ;
import csr_types        :: * ;
import Assert           :: * ;
`include "csrbox.defines"
`include "Logger.bsv"

  // Interaface declaration
  interface Ifc_csrbox_grp1;
    method Action ma_stop_count(Bit#(1) _stop);

    method Bit#(64) mv_csr_misa;
    method Bit#(32) mv_csr_mvendorid;
    method Bit#(64) mv_csr_stvec;
    method Bit#(64) mv_csr_mtvec;
    method Bit#(64) mv_csr_mstatus;
    method Bit#(64) mv_csr_marchid;
    method Bit#(64) mv_csr_mimpid;
    method Bit#(64) mv_csr_mhartid;
    method Bit#(64) mv_csr_mip;
    method Bit#(64) mv_csr_sip;
    method Bit#(64) mv_csr_mie;
    method Bit#(64) mv_csr_sie;
    method Bit#(64) mv_csr_mscratch;
    method Bit#(64) mv_csr_sscratch;
    method Bit#(64) mv_csr_sepc;
    method Bit#(64) mv_csr_stval;
    method Bit#(64) mv_csr_scause;
    method Bit#(64) mv_csr_mepc;
    method Bit#(64) mv_csr_mtval;
    method Bit#(64) mv_csr_mcause;
    method Bit#(64) mv_csr_mcycle;
    method Bit#(64) mv_csr_minstret;
    method Bit#(64) mv_csr_fcsr;
    method Bit#(64) mv_csr_time;
    method Bit#(64) mv_csr_mideleg;
    method Bit#(64) mv_csr_medeleg;
    method Bit#(64) mv_csr_pmpcfg0;
    method Bit#(30) mv_csr_pmpaddr0;
    method Bit#(30) mv_csr_pmpaddr1;
    method Bit#(30) mv_csr_pmpaddr2;
    method Bit#(30) mv_csr_pmpaddr3;
    method Bit#(32) mv_csr_mcounteren;
    method Bit#(32) mv_csr_scounteren;
    method Bit#(64) mv_csr_satp;
    method Bit#(32) mv_csr_mcountinhibit;
    method Bit#(5) mv_csr_fflags;
    method Bit#(3) mv_csr_frm;
    method Bit#(64) mv_csr_customcontrol;
    method Action ma_set_mstatus_mpie (Bit#(1) _mpie);
    method Action ma_set_mstatus_mpp (Bit#(2) _mpp);
    method Action ma_set_mstatus_mie (Bit#(1) _mie);
    method Action ma_set_mstatus_spie (Bit#(1) _spie);
    method Action ma_set_mstatus_spp (Bit#(1) _spp);
    method Action ma_set_mstatus_sie (Bit#(1) _sie);
    method Action ma_set_mstatus_upie (Bit#(1) _upie);
    method Action ma_set_mstatus_uie (Bit#(1) _uie);
    method Action ma_set_mstatus_mprv (Bit#(1) _mprv);
    method Action ma_set_mstatus_sd (Bit#(1) _sd);
    method Action ma_set_mstatus_fs (Bit#(2) _fs);
     method Action ma_set_mstatus_uxl (Bit#(2) _uxl);
    
    
    method Action ma_set_mstatus_sum (Bit#(1) _sum);
    method Action ma_set_mstatus_mxr (Bit#(1) _mxr);
    method Action ma_set_mip_meip (Bit#(1) _meip);
    method Action ma_set_mip_mtip (Bit#(1) _mtip);
    method Action ma_set_mip_msip (Bit#(1) _msip);
    method Action ma_set_mip_seip (Bit#(1) _seip);
    method Action ma_set_sepc (Bit#(64) _epc);
    method Action ma_set_stval (Bit#(64) _tval);
    method Action ma_set_scause (Bit#(64) _cause);
    method Action ma_set_mepc (Bit#(64) _mepc);
    method Action ma_set_mtval (Bit#(64) _tval);
    method Action ma_set_mcause (Bit#(64) _cause);
    method Action ma_incr_minstret(Bit#(64) incr);
    method Action ma_set_time (Bit#(64) _time);
    method Action ma_set_fflags (Bit#(5) _fflags);

    method Action ma_set_mip_debug_interrupt (Bit#(1) _debug_interrupt);    
    /*doc:method : to receive the request from the core or previous node" */
    method Action ma_core_req(CSRReq req); 

    /*doc:method : to send response to core on a hit in this node" */
    method CSRResponse mv_core_resp;

    /*doc:method: fetch from core the prvilege mode */
    method Action ma_upd_privilege (Privilege_mode prv);
    
    /*doc:method: fetch from core the virtual mode */
    method Action ma_upd_virtual (Bit#(1) _virtual);
    
    method Action ma_upd_debug_mode (Bit#(1) _dbg);
    
    /*doc:method: to forward the request to the next node on a miss in current node*/
    method ActionValue#(CSRReq) mav_fwd_req;

  endinterface

  //Module Declarations
`ifdef csrbox_grp_noinline
  (*synthesize*)
  
  (*conflict_free="ma_core_req,mv_core_resp"*)
  (*mutually_exclusive = "ma_set_mstatus_mpie, ma_core_req"*)
  (*mutually_exclusive = "ma_set_mstatus_mpp, ma_core_req"*)
  (*mutually_exclusive = "ma_set_mstatus_mie, ma_core_req"*)
  (*mutually_exclusive = "ma_set_mstatus_spie, ma_core_req"*)
  (*mutually_exclusive = "ma_set_mstatus_spp, ma_core_req"*)
  (*mutually_exclusive = "ma_set_mstatus_sie, ma_core_req"*)
  (*mutually_exclusive = "ma_set_mstatus_upie, ma_core_req"*)
  (*mutually_exclusive = "ma_set_mstatus_uie, ma_core_req"*)
  (*mutually_exclusive = "ma_set_mstatus_mprv, ma_core_req"*)
  (*mutually_exclusive = "ma_set_mstatus_sd, ma_core_req"*)
  (*mutually_exclusive = "ma_set_mstatus_fs , ma_core_req"*)
 (*mutually_exclusive = "ma_set_mstatus_uxl, ma_core_req"*)
(*mutually_exclusive="ma_set_mstatus_sum, ma_core_req"*)
(*mutually_exclusive="ma_set_mstatus_mxr ,ma_core_req"*)
  (*mutually_exclusive = "ma_set_mip_meip, ma_core_req"*)
  (*mutually_exclusive = "ma_set_mip_mtip, ma_core_req"*)
  (*mutually_exclusive = "ma_set_mip_msip, ma_core_req"*)
  (*mutually_exclusive = "ma_set_sepc, ma_core_req"*)
  (*mutually_exclusive = "ma_set_stval, ma_core_req"*)
  (*mutually_exclusive = "ma_set_scause, ma_core_req"*)
  (*mutually_exclusive = "ma_set_mepc, ma_core_req"*)
  (*mutually_exclusive = "ma_set_mtval, ma_core_req"*)
  (*mutually_exclusive = "ma_set_mcause, ma_core_req"*)
  (*preempts="ma_core_req, ma_set_fflags"*)

`endif
  module mk_csrbox_grp1(Ifc_csrbox_grp1);

    String csrbox = "";


    /*doc:wire: holds the response of this group for a csr operation request,
    for one cycle, wire is used for low latency*/
    Wire#(CSRResponse) rg_resp_to_core <- mkDWire(CSRResponse{hit:False, data:0
        `ifdef rtldump , csr_updated: False `endif });

    /*doc:fifo: fifo to forward the core request to the next group on a miss*/
    FIFOF#(CSRReq) ff_fwd_request <- mkFIFOF();

    /*doc:wire: holds the current privilege mode of the hart*/
    Wire#(Privilege_mode) wr_prv <- mkWire();
   
    /*doc:wire: holds the current state of the vs bit of the hart*/
    Wire#(Bit#(1)) wr_virtual <- mkWire();

    Wire#(Bit#(1)) wr_debug_mode <- mkWire();

    Bit#(`pmp_grain) tor = 0;
    Bit#(30) napot_mask = 0;
    Bit#(30) tor_mask = signExtend({1'b1,tor});

    Wire#(Bit#(1)) wr_ex_seip <- mkDWire(0);
    Wire#(Bit#(1)) wr_stop_count <- mkDWire(0);
    function Reg#(Bit#(26)) warlReg_misa_extensions(Reg#(Bit#(26)) r);
        return (interface Reg;
            method Bit#(26) _read = r;
            method Action _write(Bit#(26) x);
               if (True) begin
                   if (True) begin
                       let _x = x;
                       _x[25:0] = (x[25:0] & 'h14112d) | (~'h14112d & 'h0);

                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_misa_extensions

    /*doc:reg: Encodes the presence of the standard extensions, with a single bit per letter of the alphabet.*/
    Reg#(Bit#(26)) rg_misa_extensions_warl <- mkReg(1315117);
    Reg#(Bit#(26)) rg_misa_extensions = warlReg_misa_extensions(rg_misa_extensions_warl);

    function Reg#(Bit#(2)) warlReg_misa_mxl(Reg#(Bit#(2)) r);
        return (interface Reg;
            method Bit#(2) _read = r;
            method Action _write(Bit#(2) x);
               if (True) begin
                   if (( x[1:0] == 2 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_misa_mxl

    /*doc:reg: Encodes the native base integer ISA width.*/
    Reg#(Bit#(2)) rg_misa_mxl_warl <- mkReg(2);
    Reg#(Bit#(2)) rg_misa_mxl = warlReg_misa_mxl(rg_misa_mxl_warl);

    /*doc:reg: misa is a read-write register reporting the ISA supported by the hart. */
    Reg#(Bit#(64)) rg_misa = concatReg3( rg_misa_mxl , readOnlyReg(36'd0) ,rg_misa_extensions );

    /*doc:reg: 32-bit read-only register providing the JEDEC manufacturer ID of the provider of the core.*/
    Reg#(Bit#(32)) rg_mvendorid = readOnlyReg(0);

    function Reg#(Bit#(2)) warlReg_stvec_mode(Reg#(Bit#(2)) r);
        return (interface Reg;
            method Bit#(2) _read = r;
            method Action _write(Bit#(2) x);
               if (True) begin
                   if (( x[1:0] >= 0 && x[1:0] <= 1 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_stvec_mode

    /*doc:reg: Vector mode.*/
    Reg#(Bit#(2)) rg_stvec_mode_warl <- mkReg(0);
    Reg#(Bit#(2)) rg_stvec_mode = warlReg_stvec_mode(rg_stvec_mode_warl);

    function Reg#(Bit#(62)) warlReg_stvec_base(Reg#(Bit#(62)) r);
        return (interface Reg;
            method Bit#(62) _read = r;
            method Action _write(Bit#(62) x);
               if (True) begin
                   if (True) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_stvec_base

    /*doc:reg: Vector base address.*/
    Reg#(Bit#(62)) rg_stvec_base_warl <- mkReg(0);
    Reg#(Bit#(62)) rg_stvec_base = warlReg_stvec_base(rg_stvec_base_warl);

    /*doc:reg: SXLEN-bit read/write register that holds trap vector configuration. */
    Reg#(Bit#(64)) rg_stvec = concatReg2( rg_stvec_base ,rg_stvec_mode );

    function Reg#(Bit#(2)) warlReg_mtvec_mode(Reg#(Bit#(2)) r);
        return (interface Reg;
            method Bit#(2) _read = r;
            method Action _write(Bit#(2) x);
               if (True) begin
                   if (( x[1:0] >= 0 && x[1:0] <= 1 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mtvec_mode

    /*doc:reg: Vector mode.*/
    Reg#(Bit#(2)) rg_mtvec_mode_warl <- mkReg(0);
    Reg#(Bit#(2)) rg_mtvec_mode = warlReg_mtvec_mode(rg_mtvec_mode_warl);

    function Reg#(Bit#(62)) warlReg_mtvec_base(Reg#(Bit#(62)) r);
        return (interface Reg;
            method Bit#(62) _read = r;
            method Action _write(Bit#(62) x);
               if (True) begin
                   if (True) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mtvec_base

    /*doc:reg: Vector base address.*/
    Reg#(Bit#(62)) rg_mtvec_base_warl <- mkReg(0);
    Reg#(Bit#(62)) rg_mtvec_base = warlReg_mtvec_base(rg_mtvec_base_warl);

    /*doc:reg: MXLEN-bit read/write register that holds trap vector configuration. */
    Reg#(Bit#(64)) rg_mtvec = concatReg2( rg_mtvec_base ,rg_mtvec_mode );

    /*doc:reg: Stores the state of the user mode interrupts.*/
    Reg#(Bit#(1)) rg_mstatus_uie = readOnlyReg(0);

    /*doc:reg: Stores the state of the supervisor mode interrupts.*/
    Reg#(Bit#(1)) rg_mstatus_sie <- mkReg(0);

    /*doc:reg: Stores the state of the machine mode interrupts.*/
    Reg#(Bit#(1)) rg_mstatus_mie <- mkReg(0);

    /*doc:reg: Stores the state of the user mode interrupts prior to the trap.*/
    Reg#(Bit#(1)) rg_mstatus_upie = readOnlyReg(0);

    /*doc:reg: Stores the state of the supervisor mode interrupts prior to the trap.*/
    Reg#(Bit#(1)) rg_mstatus_spie <- mkReg(0);

    /*doc:reg: Stores the state of the machine mode interrupts prior to the trap.*/
    Reg#(Bit#(1)) rg_mstatus_mpie <- mkReg(0);

    /*doc:reg: Stores the previous priority mode for supervisor.*/
    Reg#(Bit#(1)) rg_mstatus_spp <- mkReg(0);

    function Reg#(Bit#(2)) warlReg_mstatus_mpp(Reg#(Bit#(2)) r);
        return (interface Reg;
            method Bit#(2) _read = r;
            method Action _write(Bit#(2) x);
               if (True) begin
                   if (( x[1:0] == 0 || x[1:0] == 1 || x[1:0] == 3 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mstatus_mpp

    /*doc:reg: Stores the previous priority mode for machine.*/
    Reg#(Bit#(2)) rg_mstatus_mpp_warl <- mkReg(0);
    Reg#(Bit#(2)) rg_mstatus_mpp = warlReg_mstatus_mpp(rg_mstatus_mpp_warl);

    function Reg#(Bit#(2)) warlReg_mstatus_fs(Reg#(Bit#(2)) r);
        return (interface Reg;
            method Bit#(2) _read = r;
            method Action _write(Bit#(2) x);
               if (True) begin
                   if (( True )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mstatus_fs

    /*doc:reg: Encodes the status of the floating-point unit, including the CSR fcsr and floating-point data registers.*/
    Reg#(Bit#(2)) rg_mstatus_fs_warl <- mkReg(0);
    Reg#(Bit#(2)) rg_mstatus_fs = warlReg_mstatus_fs(rg_mstatus_fs_warl);

    /*doc:reg: Encodes the status of additional user-mode extensions and associated state.*/
    Reg#(Bit#(2)) rg_mstatus_xs = readOnlyReg(0);

    function Reg#(Bit#(1)) warlReg_mstatus_mprv(Reg#(Bit#(1)) r);
        return (interface Reg;
            method Bit#(1) _read = r;
            method Action _write(Bit#(1) x);
               if (True) begin
                   if (( True )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mstatus_mprv

    /*doc:reg: Modifies the privilege level at which loads and stores execute in all privilege modes.*/
    Reg#(Bit#(1)) rg_mstatus_mprv_warl <- mkReg(0);
    Reg#(Bit#(1)) rg_mstatus_mprv = warlReg_mstatus_mprv(rg_mstatus_mprv_warl);

    /*doc:reg: Modifies the privilege with which S-mode loads and stores access virtual memory.*/
    Reg#(Bit#(1)) rg_mstatus_sum <- mkReg(0);

    /*doc:reg: Modifies the privilege with which loads access virtual memory.*/
    Reg#(Bit#(1)) rg_mstatus_mxr <- mkReg(0);

    /*doc:reg: Supports intercepting supervisor virtual-memory management operations.*/
    Reg#(Bit#(1)) rg_mstatus_tvm <- mkReg(0);

    /*doc:reg: Supports intercepting the WFI instruction.*/
    Reg#(Bit#(1)) rg_mstatus_tw <- mkReg(0);

    /*doc:reg: Supports intercepting the supervisor exception return instruction.*/
    Reg#(Bit#(1)) rg_mstatus_tsr <- mkReg(0);

    /*doc:reg: Controls the xlen for User mode.*/
    Reg#(Bit#(2)) rg_mstatus_uxl = readOnlyReg(2);

    /*doc:reg: Controls the value of xlen for Supervisor mode.*/
    Reg#(Bit#(2)) rg_mstatus_sxl = readOnlyReg(2);

    /*doc:reg: For any trap (access fault, page fault, or guest-page fault) that writes a guest virtual address to mtval, GVA is set to 1.*/
    Reg#(Bit#(1)) rg_mstatus_gva = readOnlyReg(0);

    /*doc:reg: Machine Previous Virtualization Mode is written by the implementation whenever a trap is taken into M-mode.*/
    Reg#(Bit#(1)) rg_mstatus_mpv = readOnlyReg(0);

    /*doc:reg: Read-only bit that summarizes whether either the FS field or XS field signals the presence of some dirty state.*/
    Reg#(Bit#(1)) rg_mstatus_sd = readOnlyReg(pack((rg_mstatus_xs == 2'b11) || (rg_mstatus_fs == 2'b11)));

    /*doc:reg: The mstatus register keeps track of and controls the hart’s current operating state. */
    Reg#(Bit#(64)) rg_mstatus = concatReg27( rg_mstatus_sd , readOnlyReg(23'd0) ,rg_mstatus_mpv ,rg_mstatus_gva , readOnlyReg(2'd0) ,rg_mstatus_sxl ,rg_mstatus_uxl , readOnlyReg(9'd0) ,rg_mstatus_tsr ,rg_mstatus_tw ,rg_mstatus_tvm ,rg_mstatus_mxr ,rg_mstatus_sum ,rg_mstatus_mprv ,rg_mstatus_xs ,rg_mstatus_fs ,rg_mstatus_mpp , readOnlyReg(2'd0) ,rg_mstatus_spp ,rg_mstatus_mpie , readOnlyReg(1'd0) ,rg_mstatus_spie ,rg_mstatus_upie ,rg_mstatus_mie , readOnlyReg(1'd0) ,rg_mstatus_sie ,rg_mstatus_uie );

    /*doc:reg: The sstatus register keeps track of the processor’s current operating state. */
    Reg#(Bit#(64)) rg_sstatus = concatReg17( rg_mstatus_sd , readOnlyReg(29'd0) ,rg_mstatus_uxl , readOnlyReg(12'd0) ,rg_mstatus_mxr ,rg_mstatus_sum , readOnlyReg(1'd0) ,rg_mstatus_xs ,rg_mstatus_fs , readOnlyReg(4'd0) ,rg_mstatus_spp , readOnlyReg(2'd0) ,rg_mstatus_spie ,rg_mstatus_upie , readOnlyReg(2'd0) ,rg_mstatus_sie ,rg_mstatus_uie );

    /*doc:reg: MXLEN-bit read-only register encoding the base microarchitecture of the hart.*/
    Reg#(Bit#(64)) rg_marchid = readOnlyReg(5);

    /*doc:reg: Provides a unique encoding of the version of the processor implementation.*/
    Reg#(Bit#(64)) rg_mimpid = readOnlyReg(0);

    /*doc:reg: MXLEN-bit read-only register containing the integer ID of the hardware thread running the code.*/
    Reg#(Bit#(64)) rg_mhartid = readOnlyReg(0);

    /*doc:reg: User Software Interrupt Pending.*/
    Reg#(Bit#(1)) rg_mip_usip = readOnlyReg(0);

    /*doc:reg: Supervisor Software Interrupt Pending.*/
    Reg#(Bit#(1)) rg_mip_ssip <- mkReg(0);

    function Reg#(Bit#(1)) warlReg_mip_vssip(Reg#(Bit#(1)) r);
        return (interface Reg;
            method Bit#(1) _read = r;
            method Action _write(Bit#(1) x);
               if (True) begin
                   if (( x[0] == 0 || x[0] == 1 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mip_vssip

    /*doc:reg: VS-level Software Interrupt Pending.*/
    Reg#(Bit#(1)) rg_mip_vssip_warl <- mkReg(0);
    Reg#(Bit#(1)) rg_mip_vssip = warlReg_mip_vssip(rg_mip_vssip_warl);

    /*doc:wire: */
    Wire#(Bit#(1)) rg_mip_msip <- mkDWire(0);

    /*doc:reg: User Timer Interrupt Pending.*/
    Reg#(Bit#(1)) rg_mip_utip = readOnlyReg(0);

    /*doc:reg: Supervisor Timer Interrupt Pending.*/
    Reg#(Bit#(1)) rg_mip_stip <- mkReg(0);

    function Reg#(Bit#(1)) warlReg_mip_vstip(Reg#(Bit#(1)) r);
        return (interface Reg;
            method Bit#(1) _read = r;
            method Action _write(Bit#(1) x);
               if (True) begin
                   if (( x[0] == 0 || x[0] == 1 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mip_vstip

    /*doc:reg: VS-level Timer Interrupt Pending.*/
    Reg#(Bit#(1)) rg_mip_vstip_warl <- mkReg(0);
    Reg#(Bit#(1)) rg_mip_vstip = warlReg_mip_vstip(rg_mip_vstip_warl);

    /*doc:wire: */
    Wire#(Bit#(1)) rg_mip_mtip <- mkDWire(0);

    /*doc:reg: User External Interrupt Pending.*/
    Reg#(Bit#(1)) rg_mip_ueip = readOnlyReg(0);

    /*doc:reg: Supervisor External Interrupt Pending.*/
    Reg#(Bit#(1)) rg_mip_seip <- mkReg(0);

    function Reg#(Bit#(1)) warlReg_mip_vseip(Reg#(Bit#(1)) r);
        return (interface Reg;
            method Bit#(1) _read = r;
            method Action _write(Bit#(1) x);
               if (True) begin
                   if (( x[0] == 0 || x[0] == 1 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mip_vseip

    /*doc:reg: VS-level External Interrupt Pending.*/
    Reg#(Bit#(1)) rg_mip_vseip_warl <- mkReg(0);
    Reg#(Bit#(1)) rg_mip_vseip = warlReg_mip_vseip(rg_mip_vseip_warl);

    /*doc:wire: */
    Wire#(Bit#(1)) rg_mip_meip <- mkDWire(0);

    /*doc:reg: HS-level External Interrupt Pending.*/
    Reg#(Bit#(1)) rg_mip_sgeip = readOnlyReg(0);

    /*doc:wire: */
    Wire#(Bit#(1)) rg_mip_debug_interrupt <- mkDWire(0);

    /*doc:reg: The mip register is an MXLEN-bit read/write register containing information on pending interrupts. */
    Reg#(Bit#(64)) rg_mip = concatReg16(  readOnlyReg(47'd0) ,readOnlyReg(rg_mip_debug_interrupt),  readOnlyReg(3'd0) ,rg_mip_sgeip ,readOnlyReg(rg_mip_meip), rg_mip_vseip ,rg_mip_seip ,rg_mip_ueip ,readOnlyReg(rg_mip_mtip), rg_mip_vstip ,rg_mip_stip ,rg_mip_utip ,readOnlyReg(rg_mip_msip), rg_mip_vssip ,rg_mip_ssip ,rg_mip_usip );

    /*doc:reg: The sip register is an SXLEN-bit read/write register containing interrupt pending bits. */
    Reg#(Bit#(64)) rg_sip = concatReg9(  readOnlyReg(54'd0) ,readOnlyReg(rg_mip_seip), rg_mip_ueip , readOnlyReg(2'd0) ,readOnlyReg(rg_mip_stip), rg_mip_utip , readOnlyReg(2'd0) ,rg_mip_ssip ,rg_mip_usip );

    /*doc:reg: User Software Interrupt enable.*/
    Reg#(Bit#(1)) rg_mie_usie = readOnlyReg(0);

    /*doc:reg: Supervisor Software Interrupt enable.*/
    Reg#(Bit#(1)) rg_mie_ssie <- mkReg(0);

    function Reg#(Bit#(1)) warlReg_mie_vssie(Reg#(Bit#(1)) r);
        return (interface Reg;
            method Bit#(1) _read = r;
            method Action _write(Bit#(1) x);
               if (True) begin
                   if (( x[0] == 0 || x[0] == 1 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mie_vssie

    /*doc:reg: VS-level Software Interrupt enable.*/
    Reg#(Bit#(1)) rg_mie_vssie_warl <- mkReg(0);
    Reg#(Bit#(1)) rg_mie_vssie = warlReg_mie_vssie(rg_mie_vssie_warl);

    /*doc:reg: Machine Software Interrupt enable.*/
    Reg#(Bit#(1)) rg_mie_msie <- mkReg(0);

    /*doc:reg: User Timer Interrupt enable.*/
    Reg#(Bit#(1)) rg_mie_utie = readOnlyReg(0);

    /*doc:reg: Supervisor Timer Interrupt enable.*/
    Reg#(Bit#(1)) rg_mie_stie <- mkReg(0);

    function Reg#(Bit#(1)) warlReg_mie_vstie(Reg#(Bit#(1)) r);
        return (interface Reg;
            method Bit#(1) _read = r;
            method Action _write(Bit#(1) x);
               if (True) begin
                   if (( x[0] == 0 || x[0] == 1 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mie_vstie

    /*doc:reg: VS-level Timer Interrupt enable.*/
    Reg#(Bit#(1)) rg_mie_vstie_warl <- mkReg(0);
    Reg#(Bit#(1)) rg_mie_vstie = warlReg_mie_vstie(rg_mie_vstie_warl);

    /*doc:reg: Machine Timer Interrupt enable.*/
    Reg#(Bit#(1)) rg_mie_mtie <- mkReg(0);

    /*doc:reg: User External Interrupt enable.*/
    Reg#(Bit#(1)) rg_mie_ueie = readOnlyReg(0);

    /*doc:reg: Supervisor External Interrupt enable.*/
    Reg#(Bit#(1)) rg_mie_seie <- mkReg(0);

    function Reg#(Bit#(1)) warlReg_mie_vseie(Reg#(Bit#(1)) r);
        return (interface Reg;
            method Bit#(1) _read = r;
            method Action _write(Bit#(1) x);
               if (True) begin
                   if (( x[0] == 0 || x[0] == 1 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mie_vseie

    /*doc:reg: VS-level External Interrupt enable.*/
    Reg#(Bit#(1)) rg_mie_vseie_warl <- mkReg(0);
    Reg#(Bit#(1)) rg_mie_vseie = warlReg_mie_vseie(rg_mie_vseie_warl);

    /*doc:reg: Machine External Interrupt enable.*/
    Reg#(Bit#(1)) rg_mie_meie <- mkReg(0);

    /*doc:reg: HS-level External Interrupt enable.*/
    Reg#(Bit#(1)) rg_mie_sgeie = readOnlyReg(0);

    /*doc:reg: */
    Reg#(Bit#(1)) rg_mie_debug_interrupt <- mkReg(1);

    /*doc:reg: The mie register is an MXLEN-bit read/write register containing interrupt enable bits. */
    Reg#(Bit#(64)) rg_mie = concatReg16(  readOnlyReg(47'd0) ,rg_mie_debug_interrupt , readOnlyReg(3'd0) ,rg_mie_sgeie ,rg_mie_meie ,rg_mie_vseie ,rg_mie_seie ,rg_mie_ueie ,rg_mie_mtie ,rg_mie_vstie ,rg_mie_stie ,rg_mie_utie ,rg_mie_msie ,rg_mie_vssie ,rg_mie_ssie ,rg_mie_usie );

    /*doc:reg: The sie register is an SXLEN-bit read/write register containing interrupt enable bits. */
    Reg#(Bit#(64)) rg_sie = concatReg9(  readOnlyReg(54'd0) ,rg_mie_seie ,rg_mie_ueie , readOnlyReg(2'd0) ,rg_mie_stie ,rg_mie_utie , readOnlyReg(2'd0) ,rg_mie_ssie ,rg_mie_usie );

    function Reg#(Bit#(64)) warlReg_mscratch(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (( True )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mscratch

    /*doc:reg: The mscratch register is an MXLEN-bit read/write register dedicated for use by machine mode.*/
    Reg#(Bit#(64)) rg_mscratch_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_mscratch = warlReg_mscratch(rg_mscratch_warl);

    function Reg#(Bit#(64)) warlReg_sscratch(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (( True )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_sscratch

    /*doc:reg: The sscratch register is an MXLEN-bit read/write register dedicated for use by machine mode.*/
    Reg#(Bit#(64)) rg_sscratch_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_sscratch = warlReg_sscratch(rg_sscratch_warl);

    function Reg#(Bit#(64)) warlReg_sepc(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (True) begin
                       let _x = x;
                       _x[63:0] = (x[63:0] & 'hfffffffffffffffe) | (~'hfffffffffffffffe & 'h0);

                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_sepc

    /*doc:reg: The sepc is a warl register that must be able to hold all valid physical and virtual addresses.*/
    Reg#(Bit#(64)) rg_sepc_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_sepc = warlReg_sepc(rg_sepc_warl);

    function Reg#(Bit#(64)) warlReg_stval(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (( True )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_stval

    /*doc:reg: The stval is a warl register that holds the address of the instruction which caused the exception.*/
    Reg#(Bit#(64)) rg_stval_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_stval = warlReg_stval(rg_stval_warl);

    function Reg#(Bit#(63)) wlrlReg_scause_exception_code(Reg#(Bit#(5)) r);
        return (interface Reg;
            method Bit#(63) _read = zeroExtend(r);
            method Action _write(Bit#(63) x);
                r._write(truncate(x));
            endmethod
        endinterface);
    endfunction: wlrlReg_scause_exception_code

    /*doc:reg: Encodes the exception code.*/
    Reg#(Bit#(5)) rg_scause_exception_code_wlrl <- mkReg(0);
    Reg#(Bit#(63)) rg_scause_exception_code = wlrlReg_scause_exception_code(rg_scause_exception_code_wlrl);

    /*doc:reg: Indicates whether the trap was due to an interrupt.*/
    Reg#(Bit#(1)) rg_scause_interrupt <- mkReg(0);

    /*doc:reg: The scause register stores the information regarding the trap. */
    Reg#(Bit#(64)) rg_scause = concatReg2( rg_scause_interrupt ,rg_scause_exception_code );

    function Reg#(Bit#(64)) warlReg_mepc(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (True) begin
                       let _x = x;
                       _x[63:0] = (x[63:0] & 'hfffffffffffffffe) | (~'hfffffffffffffffe & 'h0);

                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mepc

    /*doc:reg: The mepc is a warl register that must be able to hold all valid physical and virtual addresses.*/
    Reg#(Bit#(64)) rg_mepc_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_mepc = warlReg_mepc(rg_mepc_warl);

    function Reg#(Bit#(64)) warlReg_mtval(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (( True )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mtval

    /*doc:reg: The mtval is a warl register that holds the address of the instruction which caused the exception.*/
    Reg#(Bit#(64)) rg_mtval_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_mtval = warlReg_mtval(rg_mtval_warl);

    function Reg#(Bit#(63)) wlrlReg_mcause_exception_code(Reg#(Bit#(5)) r);
        return (interface Reg;
            method Bit#(63) _read = zeroExtend(r);
            method Action _write(Bit#(63) x);
                r._write(truncate(x));
            endmethod
        endinterface);
    endfunction: wlrlReg_mcause_exception_code

    /*doc:reg: Encodes the exception code.*/
    Reg#(Bit#(5)) rg_mcause_exception_code_wlrl <- mkReg(0);
    Reg#(Bit#(63)) rg_mcause_exception_code = wlrlReg_mcause_exception_code(rg_mcause_exception_code_wlrl);

    /*doc:reg: Indicates whether the trap was due to an interrupt.*/
    Reg#(Bit#(1)) rg_mcause_interrupt <- mkReg(0);

    /*doc:reg: The mcause register stores the information regarding the trap. */
    Reg#(Bit#(64)) rg_mcause = concatReg2( rg_mcause_interrupt ,rg_mcause_exception_code );
    Reg#(Bit#(64)) rg_mcycle[2] <- mkCReg(2,0);
    Reg#(Bit#(64)) rg_minstret[2] <- mkCReg(2,0);

    function Reg#(Bit#(5)) warlReg_fcsr_fflags(Reg#(Bit#(5)) r);
        return (interface Reg;
            method Bit#(5) _read = r;
            method Action _write(Bit#(5) x);
               if (True) begin
                   if (( True )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_fcsr_fflags

    /*doc:reg: Stores floating point accrued exceptions.*/
    Reg#(Bit#(5)) rg_fcsr_fflags_warl <- mkReg(0);
    Reg#(Bit#(5)) rg_fcsr_fflags = warlReg_fcsr_fflags(rg_fcsr_fflags_warl);

    function Reg#(Bit#(3)) warlReg_fcsr_frm(Reg#(Bit#(3)) r);
        return (interface Reg;
            method Bit#(3) _read = r;
            method Action _write(Bit#(3) x);
               if (True) begin
                   if (( True )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_fcsr_frm

    /*doc:reg: Stores Floating-Point Dynamic Rounding Mode.*/
    Reg#(Bit#(3)) rg_fcsr_frm_warl <- mkReg(0);
    Reg#(Bit#(3)) rg_fcsr_frm = warlReg_fcsr_frm(rg_fcsr_frm_warl);

    /*doc:reg: 32-bit register to hold Floating-Point Control and Status Register. */
    Reg#(Bit#(64)) rg_fcsr = concatReg3(  readOnlyReg(56'd0) ,rg_fcsr_frm ,rg_fcsr_fflags );
    Reg#(Bit#(64)) rg_time<- mkReg(0);

    function Reg#(Bit#(64)) warlReg_mideleg(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (True) begin
                       let _x = x;
                       _x[63:0] = (x[63:0] & 'hf7ff) | (~'hf7ff & 'h0);

                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mideleg

    /*doc:reg: Machine Interrupt delegation Register.*/
    Reg#(Bit#(64)) rg_mideleg_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_mideleg = warlReg_mideleg(rg_mideleg_warl);

    function Reg#(Bit#(64)) warlReg_medeleg(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (True) begin
                       let _x = x;
                       _x[63:0] = (x[63:0] & 'hf7ff) | (~'hf7ff & 'h0);

                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_medeleg

    /*doc:reg: Machine Exception delegation Register.*/
    Reg#(Bit#(64)) rg_medeleg_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_medeleg = warlReg_medeleg(rg_medeleg_warl);

    function Reg#(Bit#(8)) warlReg_pmpcfg0_pmp0cfg(Reg#(Bit#(8)) r);
        return (interface Reg;
            method Bit#(8) _read = r;
            method Action _write(Bit#(8) x);
               if( ( r[7] == 0 )  ) begin
                   if (( x[7] >= 0 && x[7] <= 1 ) && ( x[6:5] == 0 ) && ( x[4:3] != 2 ) && ( x[2:0] != 2 && x[2:0] != 6 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_pmpcfg0_pmp0cfg

    /*doc:reg: pmp configuration bits*/
    Reg#(Bit#(8)) rg_pmpcfg0_pmp0cfg_warl <- mkReg(15);
    Reg#(Bit#(8)) rg_pmpcfg0_pmp0cfg = warlReg_pmpcfg0_pmp0cfg(rg_pmpcfg0_pmp0cfg_warl);

    function Reg#(Bit#(8)) warlReg_pmpcfg0_pmp1cfg(Reg#(Bit#(8)) r);
        return (interface Reg;
            method Bit#(8) _read = r;
            method Action _write(Bit#(8) x);
               if( ( r[7] == 0 )  ) begin
                   if (( x[7] == 0 || x[7] == 1 ) && ( x[6:5] == 0 ) && ( x[4:3] != 2 ) && ( x[2:0] != 2 && x[2:0] != 6 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_pmpcfg0_pmp1cfg

    /*doc:reg: pmp configuration bits*/
    Reg#(Bit#(8)) rg_pmpcfg0_pmp1cfg_warl <- mkReg(0);
    Reg#(Bit#(8)) rg_pmpcfg0_pmp1cfg = warlReg_pmpcfg0_pmp1cfg(rg_pmpcfg0_pmp1cfg_warl);

    function Reg#(Bit#(8)) warlReg_pmpcfg0_pmp2cfg(Reg#(Bit#(8)) r);
        return (interface Reg;
            method Bit#(8) _read = r;
            method Action _write(Bit#(8) x);
               if( ( r[7] == 0 )  ) begin
                   if (( x[7] == 0 || x[7] == 1 ) && ( x[6:5] == 0 ) && ( x[4:3] != 2 ) && ( x[2:0] != 2 && x[2:0] != 6 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_pmpcfg0_pmp2cfg

    /*doc:reg: pmp configuration bits*/
    Reg#(Bit#(8)) rg_pmpcfg0_pmp2cfg_warl <- mkReg(0);
    Reg#(Bit#(8)) rg_pmpcfg0_pmp2cfg = warlReg_pmpcfg0_pmp2cfg(rg_pmpcfg0_pmp2cfg_warl);

    function Reg#(Bit#(8)) warlReg_pmpcfg0_pmp3cfg(Reg#(Bit#(8)) r);
        return (interface Reg;
            method Bit#(8) _read = r;
            method Action _write(Bit#(8) x);
               if( ( r[7] == 0 )  ) begin
                   if (( x[7] == 0 || x[7] == 1 ) && ( x[6:5] == 0 ) && ( x[4:3] != 2 ) && ( x[2:0] != 2 && x[2:0] != 6 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_pmpcfg0_pmp3cfg

    /*doc:reg: pmp configuration bits*/
    Reg#(Bit#(8)) rg_pmpcfg0_pmp3cfg_warl <- mkReg(0);
    Reg#(Bit#(8)) rg_pmpcfg0_pmp3cfg = warlReg_pmpcfg0_pmp3cfg(rg_pmpcfg0_pmp3cfg_warl);

    /*doc:reg: pmp configuration bits*/
    Reg#(Bit#(8)) rg_pmpcfg0_pmp4cfg = readOnlyReg(0);

    /*doc:reg: pmp configuration bits*/
    Reg#(Bit#(8)) rg_pmpcfg0_pmp5cfg = readOnlyReg(0);

    /*doc:reg: pmp configuration bits*/
    Reg#(Bit#(8)) rg_pmpcfg0_pmp6cfg = readOnlyReg(0);

    /*doc:reg: pmp configuration bits*/
    Reg#(Bit#(8)) rg_pmpcfg0_pmp7cfg = readOnlyReg(0);

    /*doc:reg: PMP configuration register */
    Reg#(Bit#(64)) rg_pmpcfg0 = concatReg8( rg_pmpcfg0_pmp7cfg ,rg_pmpcfg0_pmp6cfg ,rg_pmpcfg0_pmp5cfg ,rg_pmpcfg0_pmp4cfg ,rg_pmpcfg0_pmp3cfg ,rg_pmpcfg0_pmp2cfg ,rg_pmpcfg0_pmp1cfg ,rg_pmpcfg0_pmp0cfg );

    function Reg#(Bit#(30)) warlReg_pmpaddr0(Reg#(Bit#(30)) r);
        return (interface Reg;
            method Bit#(30) _read;
                if (rg_pmpcfg0_pmp0cfg[4]==1)
                    return (r | napot_mask);
                else
                    return (r & tor_mask);
            endmethod
            method Action _write(Bit#(30) x);
               if( ( rg_pmpcfg0_pmp0cfg[7] == 0 )  ) begin
                   if (True) begin
                       let _x = x;
                       _x[29:0] = (x[29:0] & 'h3ffffffe) | (~'h3ffffffe & 'h0);

                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_pmpaddr0

    /*doc:reg: Physical memory protection address register*/
    Reg#(Bit#(30)) rg_pmpaddr0_warl <- mkReg(1073741822);
    Reg#(Bit#(30)) rg_pmpaddr0 = warlReg_pmpaddr0(rg_pmpaddr0_warl);

    function Reg#(Bit#(30)) warlReg_pmpaddr1(Reg#(Bit#(30)) r);
        return (interface Reg;
            method Bit#(30) _read;
                if (rg_pmpcfg0_pmp1cfg[4]==1)
                    return (r | napot_mask);
                else
                    return (r & tor_mask);
            endmethod
            method Action _write(Bit#(30) x);
               if( ( rg_pmpcfg0_pmp1cfg[7] == 0 )  ) begin
                   if (True) begin
                       let _x = x;
                       _x[29:0] = (x[29:0] & 'h3ffffffe) | (~'h3ffffffe & 'h0);

                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_pmpaddr1

    /*doc:reg: Physical memory protection address register*/
    Reg#(Bit#(30)) rg_pmpaddr1_warl <- mkReg(0);
    Reg#(Bit#(30)) rg_pmpaddr1 = warlReg_pmpaddr1(rg_pmpaddr1_warl);

    function Reg#(Bit#(30)) warlReg_pmpaddr2(Reg#(Bit#(30)) r);
        return (interface Reg;
            method Bit#(30) _read;
                if (rg_pmpcfg0_pmp2cfg[4]==1)
                    return (r | napot_mask);
                else
                    return (r & tor_mask);
            endmethod
            method Action _write(Bit#(30) x);
               if( ( rg_pmpcfg0_pmp2cfg[7] == 0 )  ) begin
                   if (True) begin
                       let _x = x;
                       _x[29:0] = (x[29:0] & 'h3ffffffe) | (~'h3ffffffe & 'h0);

                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_pmpaddr2

    /*doc:reg: Physical memory protection address register*/
    Reg#(Bit#(30)) rg_pmpaddr2_warl <- mkReg(0);
    Reg#(Bit#(30)) rg_pmpaddr2 = warlReg_pmpaddr2(rg_pmpaddr2_warl);

    function Reg#(Bit#(30)) warlReg_pmpaddr3(Reg#(Bit#(30)) r);
        return (interface Reg;
            method Bit#(30) _read;
                if (rg_pmpcfg0_pmp3cfg[4]==1)
                    return (r | napot_mask);
                else
                    return (r & tor_mask);
            endmethod
            method Action _write(Bit#(30) x);
               if( ( rg_pmpcfg0_pmp3cfg[7] == 0 )  ) begin
                   if (True) begin
                       let _x = x;
                       _x[29:0] = (x[29:0] & 'h3ffffffe) | (~'h3ffffffe & 'h0);

                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_pmpaddr3

    /*doc:reg: Physical memory protection address register*/
    Reg#(Bit#(30)) rg_pmpaddr3_warl <- mkReg(0);
    Reg#(Bit#(30)) rg_pmpaddr3 = warlReg_pmpaddr3(rg_pmpaddr3_warl);

    function Reg#(Bit#(32)) warlReg_mcounteren(Reg#(Bit#(32)) r);
        return (interface Reg;
            method Bit#(32) _read = r;
            method Action _write(Bit#(32) x);
               if (True) begin
                   if (True) begin
                       let _x = x;
                       _x[31:0] = (x[31:0] & 'h1f) | (~'h1f & 'h0);

                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mcounteren

    /*doc:reg: The mcounteren is a 32-bit register that controls the availability of the hardware performance-monitoring counters to the next-lowest privileged mode.*/
    Reg#(Bit#(32)) rg_mcounteren_warl <- mkReg(0);
    Reg#(Bit#(32)) rg_mcounteren = warlReg_mcounteren(rg_mcounteren_warl);

    function Reg#(Bit#(32)) warlReg_scounteren(Reg#(Bit#(32)) r);
        return (interface Reg;
            method Bit#(32) _read = r;
            method Action _write(Bit#(32) x);
               if (True) begin
                   if (True) begin
                       let _x = x;
                       _x[31:0] = (x[31:0] & 'h1f) | (~'h1f & 'h0);

                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_scounteren

    /*doc:reg: The scounteren is a 32-bit register that controls the availability of the hardware performance-monitoring counters to the next-lowest privileged mode.*/
    Reg#(Bit#(32)) rg_scounteren_warl <- mkReg(0);
    Reg#(Bit#(32)) rg_scounteren = warlReg_scounteren(rg_scounteren_warl);

    function Reg#(Bit#(44)) warlReg_satp_ppn(Reg#(Bit#(44)) r);
        return (interface Reg;
            method Bit#(44) _read = r;
            method Action _write(Bit#(44) x);
               if (True) begin
                   if (( True )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_satp_ppn

    /*doc:reg: Physical Page Number*/
    Reg#(Bit#(44)) rg_satp_ppn_warl <- mkReg(0);
    Reg#(Bit#(44)) rg_satp_ppn = warlReg_satp_ppn(rg_satp_ppn_warl);

    function Reg#(Bit#(16)) warlReg_satp_asid(Reg#(Bit#(16)) r);
        return (interface Reg;
            method Bit#(16) _read = r;
            method Action _write(Bit#(16) x);
               if (True) begin
                   if (( x[15:0] >= 0 && x[15:0] <= 255 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_satp_asid

    /*doc:reg: Address Space identifier.*/
    Reg#(Bit#(16)) rg_satp_asid_warl <- mkReg(0);
    Reg#(Bit#(16)) rg_satp_asid = warlReg_satp_asid(rg_satp_asid_warl);

    function Reg#(Bit#(4)) warlReg_satp_mode(Reg#(Bit#(4)) r);
        return (interface Reg;
            method Bit#(4) _read = r;
            method Action _write(Bit#(4) x);
               if (True) begin
                   if (( x[3:0] == 0 || x[3:0] == 8 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_satp_mode

    /*doc:reg: Vector mode.*/
    Reg#(Bit#(4)) rg_satp_mode_warl <- mkReg(0);
    Reg#(Bit#(4)) rg_satp_mode = warlReg_satp_mode(rg_satp_mode_warl);

    /*doc:reg: SXLEN-bit register which controls supervisor-mode address translation and protection */
    Reg#(Bit#(64)) rg_satp = concatReg3( rg_satp_mode ,rg_satp_asid ,rg_satp_ppn );

    /*doc:reg: The mcountinhibit is a 32-bit WARL register that controls which of the hardware performance-monitoring counters increment.*/
    Reg#(Bit#(32)) rg_mcountinhibit = readOnlyReg(0);

    /*doc:reg: bit for cache-enable of instruction cache, part of rg_customcontrol*/
    Reg#(Bit#(1)) rg_customcontrol_ienable = readOnlyReg(1);

    /*doc:reg: bit for cache-enable of data cache, part of rg_customcontrol*/
    Reg#(Bit#(1)) rg_customcontrol_denable = readOnlyReg(1);

    /*doc:reg: bit for enabling branch predictor unit, part of rg_customcontrol*/
    Reg#(Bit#(1)) rg_customcontrol_bpuenable = readOnlyReg(1);

    /*doc:reg: bit for enabling arithmetic exceptions, part of rg_customcontrol*/
    Reg#(Bit#(1)) rg_customcontrol_arith_excep = readOnlyReg(0);

    /*doc:reg: bit for enabling debugger on the current hart*/
    Reg#(Bit#(1)) rg_customcontrol_debug_enable = readOnlyReg(1);

    /*doc:reg: the register holds enable bits for arithmetic exceptions, branch predictor unit, i-cache, d-cache units */
    Reg#(Bit#(64)) rg_customcontrol = concatReg6(  readOnlyReg(59'd0) ,rg_customcontrol_debug_enable ,rg_customcontrol_arith_excep ,rg_customcontrol_bpuenable ,rg_customcontrol_denable ,rg_customcontrol_ienable );
    rule rl_increment_cycle;
      if (wr_stop_count == 0 )
        rg_mcycle[0] <= rg_mcycle[0] + 1;
    endrule
 
    method Action ma_core_req(CSRReq req);
        `logLevel( csrbox_grp1, 1, $format("csrbox_grp1: received req: ", fshow(req)))
        Bit#(2) op = req.funct3; 
        case (req.csr_address)             `MISA:begin
              Bit#(64) readdata = zeroExtend(rg_misa);
              let word = fn_csr_op(req.writedata, readdata, op);
              word[3] = word[3] & word[5]; // is D is being disabled, then disable F as well.
              Bool supress_changes = rg_misa[2]== 1 && word[2]==0 && req.pc_1 == 1;
              if (!supress_changes)
                rg_misa <= truncate(word);
              rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump, csr_updated: !supress_changes `endif };
            end

            `MVENDORID : begin
                Bit#(64) readdata = zeroExtend(rg_mvendorid);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump , csr_updated : False `endif };
            end

            `STVEC : begin
                Bit#(64) readdata = zeroExtend(rg_stvec);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_stvec <= truncate(word);
            end

            `MTVEC : begin
                Bit#(64) readdata = zeroExtend(rg_mtvec);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_mtvec <= truncate(word);
            end

            `MSTATUS : begin
                Bit#(64) readdata = zeroExtend(rg_mstatus);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_mstatus <= truncate(word);
            end

            `SSTATUS : begin
                Bit#(64) readdata = zeroExtend(rg_sstatus);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_sstatus <= truncate(word);
            end

            `MARCHID : begin
                Bit#(64) readdata = zeroExtend(rg_marchid);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump , csr_updated : False `endif };
            end

            `MIMPID : begin
                Bit#(64) readdata = zeroExtend(rg_mimpid);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump , csr_updated : False `endif };
            end

            `MHARTID : begin
                Bit#(64) readdata = zeroExtend(rg_mhartid);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump , csr_updated : False `endif };
            end
            `MIP:begin
                Bit#(64) readdata = truncate(rg_mip);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata | {'d0,wr_ex_seip,9'd0} `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, truncate(rg_mip), op);
                rg_mip <= word;
            end
            `SIP : begin
                Bit#(64) readdata = truncate(rg_sip);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata | {'d0,wr_ex_seip,9'd0}  `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, truncate(rg_sip), op);
                rg_sip <= word;
            end

            `MIE : begin
                Bit#(64) readdata = zeroExtend(rg_mie);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_mie <= truncate(word);
            end

            `SIE : begin
                Bit#(64) readdata = zeroExtend(rg_sie);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_sie <= truncate(word);
            end

            `MSCRATCH : begin
                Bit#(64) readdata = zeroExtend(rg_mscratch);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_mscratch <= truncate(word);
            end

            `SSCRATCH : begin
                Bit#(64) readdata = zeroExtend(rg_sscratch);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_sscratch <= truncate(word);
            end

            `SEPC : begin
                Bit#(64) readdata = zeroExtend(rg_sepc);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_sepc <= truncate(word);
            end

            `STVAL : begin
                Bit#(64) readdata = zeroExtend(rg_stval);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_stval <= truncate(word);
            end

            `SCAUSE : begin
                Bit#(64) readdata = zeroExtend(rg_scause);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_scause <= truncate(word);
            end

            `MEPC : begin
                Bit#(64) readdata = zeroExtend(rg_mepc);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_mepc <= truncate(word);
            end

            `MTVAL : begin
                Bit#(64) readdata = zeroExtend(rg_mtval);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_mtval <= truncate(word);
            end

            `MCAUSE : begin
                Bit#(64) readdata = zeroExtend(rg_mcause);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_mcause <= truncate(word);
            end
            `MCYCLE : begin
                Bit#(64) readdata = truncate(rg_mcycle[1]);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                rg_mcycle[1][64-1:0] <= word;
            end
            `MINSTRET : begin
                Bit#(64) readdata = truncate(rg_minstret[0]);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                rg_minstret[0][64-1:0] <= word;
            end
            `FCSR: begin
                Bit#(64) readdata = zeroExtend(rg_fcsr);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                rg_fcsr <= word;
                rg_mstatus_fs <= 2'b11;
            end
            `TIME : begin
                Bit#(64) readdata = truncate(rg_time);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump ,csr_updated: True `endif };
            end
            `MIDELEG : begin
                        Bit#(64) readdata = zeroExtend(rg_mideleg);
                        rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump ,csr_updated: True `endif };
                        let word = fn_csr_op(req.writedata, readdata, op);
                        word[10]= word[10] | rg_misa[7] ;
                        word[6]= word[6] | rg_misa[7] ;
                        word[2]= word[2] | rg_misa[7] ;
                         rg_mideleg <= truncate(word);
                    end

            `MEDELEG : begin
                Bit#(64) readdata = zeroExtend(rg_medeleg);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_medeleg <= truncate(word);
            end

            `PMPCFG0 : begin
                Bit#(64) readdata = zeroExtend(rg_pmpcfg0);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_pmpcfg0 <= truncate(word);
            end

            `PMPADDR0 : begin
                Bit#(64) readdata = zeroExtend(rg_pmpaddr0);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_pmpaddr0 <= truncate(word);
            end

            `PMPADDR1 : begin
                Bit#(64) readdata = zeroExtend(rg_pmpaddr1);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_pmpaddr1 <= truncate(word);
            end

            `PMPADDR2 : begin
                Bit#(64) readdata = zeroExtend(rg_pmpaddr2);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_pmpaddr2 <= truncate(word);
            end

            `PMPADDR3 : begin
                Bit#(64) readdata = zeroExtend(rg_pmpaddr3);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_pmpaddr3 <= truncate(word);
            end

            `MCOUNTEREN : begin
                Bit#(64) readdata = zeroExtend(rg_mcounteren);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_mcounteren <= truncate(word);
            end

            `SCOUNTEREN : begin
                Bit#(64) readdata = zeroExtend(rg_scounteren);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_scounteren <= truncate(word);
            end
            `SATP : begin
                Bit#(64) readdata = zeroExtend(rg_satp);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                if (word[63:60] == 0||word[63:60] == 8)
                  rg_satp <= truncate(word);
            end

            `MCOUNTINHIBIT : begin
                Bit#(64) readdata = zeroExtend(rg_mcountinhibit);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_mcountinhibit <= truncate(word);
            end
            `FFLAGS: begin
                Bit#(64) readdata = zeroExtend(rg_fcsr_fflags);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                rg_fcsr_fflags <= truncate(word);
                rg_mstatus_fs <= 2'b11;
            end
            `FRM: begin
              Bit#(64) readdata = zeroExtend(rg_fcsr_frm);
              rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump ,csr_updated: True `endif };
              let word = fn_csr_op(req.writedata, readdata, op);
              rg_fcsr_frm <= truncate(word);
              rg_mstatus_fs <= 2'b11;
            end
            `CYCLE : begin
                Bit#(64) readdata = truncate(rg_mcycle[1]);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump ,csr_updated: True `endif };
            end
            `INSTRET : begin
                Bit#(64) readdata = truncate(rg_minstret[0]);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump ,csr_updated: True `endif };
            end

            `CUSTOMCONTROL : begin
                Bit#(64) readdata = zeroExtend(rg_customcontrol);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_customcontrol <= truncate(word);
            end

            default: begin
                ff_fwd_request.enq(req);
                `logLevel( csrbox_grp1, 1, $format("csrbox_grp1: fwding req to next group"))
                rg_resp_to_core <= CSRResponse{hit: False, data: 0 `ifdef rtldump , csr_updated : False `endif };
            end
        endcase
        endmethod
    
    method mv_csr_misa = rg_misa;

    method mv_csr_mvendorid = rg_mvendorid;

    method mv_csr_stvec = rg_stvec;

    method mv_csr_mtvec = rg_mtvec;

    method mv_csr_mstatus = rg_mstatus;

    method mv_csr_marchid = rg_marchid;

    method mv_csr_mimpid = rg_mimpid;

    method mv_csr_mhartid = rg_mhartid;

    method mv_csr_mip = rg_mip | {'d0,wr_ex_seip,9'd0};

    method mv_csr_sip = rg_sip | {'d0,wr_ex_seip,9'd0};

    method mv_csr_mie = rg_mie;

    method mv_csr_sie = rg_sie;

    method mv_csr_mscratch = rg_mscratch;

    method mv_csr_sscratch = rg_sscratch;

    method mv_csr_sepc = rg_sepc;

    method mv_csr_stval = rg_stval;

    method mv_csr_scause = rg_scause;

    method mv_csr_mepc = rg_mepc;

    method mv_csr_mtval = rg_mtval;

    method mv_csr_mcause = rg_mcause;

    method mv_csr_mcycle = truncate(rg_mcycle[1]);

    method mv_csr_minstret = truncate(rg_minstret[1]);

    method mv_csr_fcsr = rg_fcsr;

    method mv_csr_time = truncate(rg_time);

    method mv_csr_mideleg = rg_mideleg;

    method mv_csr_medeleg = rg_medeleg;

    method mv_csr_pmpcfg0 = rg_pmpcfg0;

    method mv_csr_pmpaddr0 = rg_pmpaddr0;

    method mv_csr_pmpaddr1 = rg_pmpaddr1;

    method mv_csr_pmpaddr2 = rg_pmpaddr2;

    method mv_csr_pmpaddr3 = rg_pmpaddr3;

    method mv_csr_mcounteren = rg_mcounteren;

    method mv_csr_scounteren = rg_scounteren;

    method mv_csr_satp = rg_satp;

    method mv_csr_mcountinhibit = rg_mcountinhibit;

    method mv_csr_fflags = rg_fcsr_fflags;

    method mv_csr_frm = rg_fcsr_frm;

    method mv_csr_customcontrol = rg_customcontrol;
    method Action ma_set_mstatus_mpie (Bit#(1) _mpie); rg_mstatus_mpie <= _mpie; endmethod
    method Action ma_set_mstatus_mpp (Bit#(2) _mpp); rg_mstatus_mpp <= _mpp; endmethod 
    method Action ma_set_mstatus_mie (Bit#(1) _mie); rg_mstatus_mie <= _mie; endmethod
    method Action ma_set_mstatus_spie (Bit#(1) _spie); rg_mstatus_spie <= _spie; endmethod
    method Action ma_set_mstatus_spp (Bit#(1) _spp); rg_mstatus_spp <= _spp; endmethod
    method Action ma_set_mstatus_sie (Bit#(1) _sie); rg_mstatus_sie <= _sie; endmethod
    method Action ma_set_mstatus_upie (Bit#(1) _upie); rg_mstatus_upie <= _upie; endmethod
    method Action ma_set_mstatus_uie (Bit#(1) _uie); rg_mstatus_uie <= _uie; endmethod
    method Action ma_set_mstatus_mprv (Bit#(1) _mprv); rg_mstatus_mprv <= _mprv; endmethod
    method Action ma_set_mstatus_fs (Bit#(2) _fs); rg_mstatus_fs <= _fs; endmethod
     method Action ma_set_mstatus_uxl (Bit#(2) _uxl); rg_mstatus_uxl <= _uxl; endmethod
    method Action ma_set_mstatus_sum (Bit#(1) _sum); rg_mstatus_sum <= _sum; endmethod
    method Action ma_set_mstatus_mxr (Bit#(1) _mxr); rg_mstatus_mxr <= _mxr; endmethod
    method Action ma_set_mstatus_sd (Bit#(1) _sd); rg_mstatus_sd <= _sd; endmethod


    method Action ma_set_mip_meip (Bit#(1) _meip);
      rg_mip_meip <= _meip;
    endmethod
    method Action ma_set_mip_mtip (Bit#(1) _mtip);
      rg_mip_mtip <= _mtip;
    endmethod
    method Action ma_set_mip_msip (Bit#(1) _msip);
      rg_mip_msip <= _msip;
    endmethod
    method Action ma_set_mip_seip (Bit#(1) _seip);
      wr_ex_seip <= _seip;
    endmethod
    method Action ma_set_sepc (Bit#(64) _epc);
      rg_sepc <= _epc;
    endmethod
    method Action ma_set_stval (Bit#(64) _tval);
      rg_stval <= _tval;
    endmethod
    method Action ma_set_scause (Bit#(64) _cause);
      rg_scause <= _cause;
    endmethod
    method Action ma_set_mepc (Bit#(64) _mepc);
      rg_mepc <= _mepc;
    endmethod
    method Action ma_set_mtval (Bit#(64) _tval);
      rg_mtval <= _tval;
    endmethod
    method Action ma_set_mcause (Bit#(64) _cause);
      rg_mcause <= _cause;
    endmethod
    method Action ma_incr_minstret(Bit#(64) incr);
      if (wr_stop_count == 0)
        rg_minstret[1] <= rg_minstret[1] + incr;
    endmethod
    method Action ma_set_time (Bit#(64) _time);
      rg_time <= _time;
    endmethod
    method Action ma_set_fflags (Bit#(5) _fflags);
      if((_fflags|truncate(rg_fcsr_fflags)) != truncate(rg_fcsr_fflags))begin
        rg_fcsr_fflags <= zeroExtend(_fflags|truncate(rg_fcsr_fflags));
        rg_mstatus_fs <= 'b11;
      end
    endmethod
    method Action ma_stop_count(Bit#(1) _stop);
      wr_stop_count <= _stop;
    endmethod

    method Action ma_set_mip_debug_interrupt (Bit#(1) _debug_interrupt);
        rg_mip_debug_interrupt <= _debug_interrupt;
    endmethod:ma_set_mip_debug_interrupt

    method mv_core_resp = rg_resp_to_core;

    method Action ma_upd_privilege (Privilege_mode prv);
        wr_prv <= prv;
    endmethod
    
    method Action ma_upd_virtual (Bit#(1) _virtual);
         wr_virtual <= _virtual;
    endmethod
    method Action ma_upd_debug_mode (Bit#(1) _dbg);
        wr_debug_mode <= _dbg;
    endmethod
        method ActionValue#(CSRReq) mav_fwd_req;
            ff_fwd_request.deq;
            return ff_fwd_request.first();
        endmethod

  endmodule 
endpackage 
